
package alu_pkg;

    `include "alu_sequence_item.sv"
    `include "alu_sequence.sv"
    `include "alu_sequencer.sv"
    `include "alu_driver.sv"
    `include "alu_a_monitor.sv"
    `include "alu_p_monitor.sv"
    `include "alu_agent.sv"
    `include "alu_scoreboard.sv"
    `include "alu_env.sv"
    `include "alu_test.sv"
    
endpackage: alu_pkg
